/************************************************************************************
 * Ask me anything: via repo/issue, or e-mail: vencifreeman16@sjtu.edu.cn.          *
 * Author: @VenciFreeman (GitHub), copyright 2019.									*
 * School: Shanghai Jiao Tong University.											*
 * Description:                                                                     *
 * Do some operations according to ALUop and the 2 source oprands.					*
 * Details:                                                                         *
 * - Use the ALUop and the two source operands decoded in id.v to perform the 		*
 *   corresponding operation;                                                       *
 * - If ALUop indicates that it's an addition operation, the two operands will be 	*
 *	 added;																			*
 * - The sub operation can be implemented by complement, etc.		                *
 * History:																			*
 * - 19/12/05: Create this file.													*
 * Notes:																			*
 ************************************************************************************/

module ex(
	
	input wire rst,
	input wire	   ALUop,
	input wire	   _srcop1_,
	input wire	   _srcop2_,
	output wire	   _output_

);	

always @ (*) begin

end	

endmodule